module app(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h0c001403;
30'h00000002: inst = 32'h37bdf000;
30'h00000003: inst = 32'h27bdffc8;
30'h00000004: inst = 32'hafbf0034;
30'h00000005: inst = 32'hafb00028;
30'h00000006: inst = 32'hafb1002c;
30'h00000007: inst = 32'hafa00020;
30'h00000008: inst = 32'h3c028000;
30'h00000009: inst = 32'h34420050;
30'h0000000a: inst = 32'h8c420000;
30'h0000000b: inst = 32'h00000000;
30'h0000000c: inst = 32'h30420001;
30'h0000000d: inst = 32'h14400005;
30'h0000000e: inst = 32'h00000000;
30'h0000000f: inst = 32'h00000000;
30'h00000010: inst = 32'h00000000;
30'h00000011: inst = 32'h08001408;
30'h00000012: inst = 32'h00000000;
30'h00000013: inst = 32'h3c028000;
30'h00000014: inst = 32'h34420050;
30'h00000015: inst = 32'h8c420000;
30'h00000016: inst = 32'h00000000;
30'h00000017: inst = 32'h30420001;
30'h00000018: inst = 32'h10400005;
30'h00000019: inst = 32'h00000000;
30'h0000001a: inst = 32'h00000000;
30'h0000001b: inst = 32'h00000000;
30'h0000001c: inst = 32'h08001413;
30'h0000001d: inst = 32'h00000000;
30'h0000001e: inst = 32'h3c028000;
30'h0000001f: inst = 32'h34420050;
30'h00000020: inst = 32'h8c420000;
30'h00000021: inst = 32'h00000000;
30'h00000022: inst = 32'h30420001;
30'h00000023: inst = 32'hafa20024;
30'h00000024: inst = 32'h3c028000;
30'h00000025: inst = 32'h34420050;
30'h00000026: inst = 32'h8c420000;
30'h00000027: inst = 32'h00000000;
30'h00000028: inst = 32'h30420001;
30'h00000029: inst = 32'h1440000f;
30'h0000002a: inst = 32'h00000000;
30'h0000002b: inst = 32'h3c021001;
30'h0000002c: inst = 32'h3c031000;
30'h0000002d: inst = 32'h34500000;
30'h0000002e: inst = 32'h24715298;
30'h0000002f: inst = 32'hae300000;
30'h00000030: inst = 32'h3404ff00;
30'h00000031: inst = 32'h0c001457;
30'h00000032: inst = 32'h00000000;
30'h00000033: inst = 32'h3c028000;
30'h00000034: inst = 32'h8e230000;
30'h00000035: inst = 32'h00000000;
30'h00000036: inst = 32'h3c041040;
30'h00000037: inst = 32'h08001446;
30'h00000038: inst = 32'h00000000;
30'h00000039: inst = 32'h3c021001;
30'h0000003a: inst = 32'h3c031000;
30'h0000003b: inst = 32'h34500000;
30'h0000003c: inst = 32'h24715298;
30'h0000003d: inst = 32'hae300000;
30'h0000003e: inst = 32'h3c0200ff;
30'h0000003f: inst = 32'h3444ffff;
30'h00000040: inst = 32'h0c001457;
30'h00000041: inst = 32'h00000000;
30'h00000042: inst = 32'h3c028000;
30'h00000043: inst = 32'h8e230000;
30'h00000044: inst = 32'h00000000;
30'h00000045: inst = 32'h3c041080;
30'h00000046: inst = 32'h34840000;
30'h00000047: inst = 32'h34450040;
30'h00000048: inst = 32'hac600000;
30'h00000049: inst = 32'h34420030;
30'h0000004a: inst = 32'haca40000;
30'h0000004b: inst = 32'hac500000;
30'h0000004c: inst = 32'h3c028000;
30'h0000004d: inst = 32'h8fa30024;
30'h0000004e: inst = 32'h00000000;
30'h0000004f: inst = 32'h34420050;
30'h00000050: inst = 32'h8c420000;
30'h00000051: inst = 32'h00000000;
30'h00000052: inst = 32'h30420001;
30'h00000053: inst = 32'h1062fff8;
30'h00000054: inst = 32'h00000000;
30'h00000055: inst = 32'h0800141e;
30'h00000056: inst = 32'h00000000;
30'h00000057: inst = 32'h27bdffe8;
30'h00000058: inst = 32'h3c021000;
30'h00000059: inst = 32'h3c030100;
30'h0000005a: inst = 32'h34630000;
30'h0000005b: inst = 32'h24425298;
30'h0000005c: inst = 32'hafa40010;
30'h0000005d: inst = 32'h00831821;
30'h0000005e: inst = 32'h8c440000;
30'h0000005f: inst = 32'h00000000;
30'h00000060: inst = 32'hac830000;
30'h00000061: inst = 32'h8c430000;
30'h00000062: inst = 32'h00000000;
30'h00000063: inst = 32'h24630004;
30'h00000064: inst = 32'hac430000;
30'h00000065: inst = 32'h27bd0018;
30'h00000066: inst = 32'h03e00008;
30'h00000067: inst = 32'h00000000;
30'h00000068: inst = 32'h27bdffd8;
30'h00000069: inst = 32'hafa40014;
30'h0000006a: inst = 32'hafa50018;
30'h0000006b: inst = 32'hafa6001c;
30'h0000006c: inst = 32'h8fa20038;
30'h0000006d: inst = 32'h00000000;
30'h0000006e: inst = 32'hafa70020;
30'h0000006f: inst = 32'hafa20024;
30'h00000070: inst = 32'h27bd0028;
30'h00000071: inst = 32'h03e00008;
30'h00000072: inst = 32'h00000000;
30'h00000073: inst = 32'h27bdffe0;
30'h00000074: inst = 32'hafa40010;
30'h00000075: inst = 32'hafa50014;
30'h00000076: inst = 32'hafa00018;
30'h00000077: inst = 32'h8fa20014;
30'h00000078: inst = 32'h00000000;
30'h00000079: inst = 32'h8fa30010;
30'h0000007a: inst = 32'h00000000;
30'h0000007b: inst = 32'h0043102a;
30'h0000007c: inst = 32'h1040000d;
30'h0000007d: inst = 32'h00000000;
30'h0000007e: inst = 32'h8fa20018;
30'h0000007f: inst = 32'h00000000;
30'h00000080: inst = 32'h24420001;
30'h00000081: inst = 32'hafa20018;
30'h00000082: inst = 32'h8fa20010;
30'h00000083: inst = 32'h00000000;
30'h00000084: inst = 32'h8fa30014;
30'h00000085: inst = 32'h00000000;
30'h00000086: inst = 32'h00431023;
30'h00000087: inst = 32'hafa20010;
30'h00000088: inst = 32'h08001477;
30'h00000089: inst = 32'h00000000;
30'h0000008a: inst = 32'h8fa20018;
30'h0000008b: inst = 32'h00000000;
30'h0000008c: inst = 32'h27bd0020;
30'h0000008d: inst = 32'h03e00008;
30'h0000008e: inst = 32'h00000000;
30'h0000008f: inst = 32'h27bdffe8;
30'h00000090: inst = 32'hafa40010;
30'h00000091: inst = 32'hafa50014;
30'h00000092: inst = 32'h8fa20010;
30'h00000093: inst = 32'h00000000;
30'h00000094: inst = 32'h8fa30014;
30'h00000095: inst = 32'h00000000;
30'h00000096: inst = 32'h0043102a;
30'h00000097: inst = 32'h14400009;
30'h00000098: inst = 32'h00000000;
30'h00000099: inst = 32'h8fa20010;
30'h0000009a: inst = 32'h00000000;
30'h0000009b: inst = 32'h8fa30014;
30'h0000009c: inst = 32'h00000000;
30'h0000009d: inst = 32'h00431023;
30'h0000009e: inst = 32'hafa20010;
30'h0000009f: inst = 32'h08001492;
30'h000000a0: inst = 32'h00000000;
30'h000000a1: inst = 32'h8fa20010;
30'h000000a2: inst = 32'h00000000;
30'h000000a3: inst = 32'h27bd0018;
30'h000000a4: inst = 32'h03e00008;
30'h000000a5: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
