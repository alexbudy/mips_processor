module isr(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h401a6800;
30'h00000001: inst = 32'h401b6000;
30'h00000002: inst = 32'h00000000;
30'h00000003: inst = 32'h337bfc00;
30'h00000004: inst = 32'h035bd024;
30'h00000005: inst = 32'h335b8000;
30'h00000006: inst = 32'h17600003;
30'h00000007: inst = 32'h00000000;
30'h00000008: inst = 32'h0800002d;
30'h00000009: inst = 32'h00000000;
30'h0000000a: inst = 32'h401b5800;
30'h0000000b: inst = 32'h241a000a;
30'h0000000c: inst = 32'h035bd021;
30'h0000000d: inst = 32'h409a5800;
30'h0000000e: inst = 32'h3c1a1000;
30'h0000000f: inst = 32'h375a00b0;
30'h00000010: inst = 32'h8f5b0000;
30'h00000011: inst = 32'h00000000;
30'h00000012: inst = 32'h277b0001;
30'h00000013: inst = 32'haf5b0000;
30'h00000014: inst = 32'h241a003c;
30'h00000015: inst = 32'h175b000c;
30'h00000016: inst = 32'h00000000;
30'h00000017: inst = 32'h0000d821;
30'h00000018: inst = 32'h3c1a1000;
30'h00000019: inst = 32'h375a00b0;
30'h0000001a: inst = 32'haf5b0000;
30'h0000001b: inst = 32'h3c1a1000;
30'h0000001c: inst = 32'h375a00b4;
30'h0000001d: inst = 32'h8f5b0000;
30'h0000001e: inst = 32'h00000000;
30'h0000001f: inst = 32'h277b0001;
30'h00000020: inst = 32'h08000022;
30'h00000021: inst = 32'haf5b0000;
30'h00000022: inst = 32'h3c1a1000;
30'h00000023: inst = 32'h375a00c8;
30'h00000024: inst = 32'h8f5b0000;
30'h00000025: inst = 32'h241a0001;
30'h00000026: inst = 32'h175b0006;
30'h00000027: inst = 32'h00000000;
30'h00000028: inst = 32'h241a004d;
30'h00000029: inst = 32'h3c1b8000;
30'h0000002a: inst = 32'h377b0008;
30'h0000002b: inst = 32'h0800002d;
30'h0000002c: inst = 32'haf7a0000;
30'h0000002d: inst = 32'h401b6000;
30'h0000002e: inst = 32'h00000000;
30'h0000002f: inst = 32'h377b0001;
30'h00000030: inst = 32'h401a7000;
30'h00000031: inst = 32'h409b6000;
30'h00000032: inst = 32'h03400008;
30'h00000033: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
