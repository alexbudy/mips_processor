module app(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h3c1d1000;
30'h00000001: inst = 32'h0c001403;
30'h00000002: inst = 32'h37bd7000;
30'h00000003: inst = 32'h27bdffd8;
30'h00000004: inst = 32'hafa00010;
30'h00000005: inst = 32'hafa00014;
30'h00000006: inst = 32'h3c0200ff;
30'h00000007: inst = 32'hafa00018;
30'h00000008: inst = 32'h3442ffff;
30'h00000009: inst = 32'hafa0001c;
30'h0000000a: inst = 32'hafa20020;
30'h0000000b: inst = 32'hafa00024;
30'h0000000c: inst = 32'h3c020009;
30'h0000000d: inst = 32'h34425e6f;
30'h0000000e: inst = 32'h8fa30024;
30'h0000000f: inst = 32'h00000000;
30'h00000010: inst = 32'h0043102a;
30'h00000011: inst = 32'h14400010;
30'h00000012: inst = 32'h00000000;
30'h00000013: inst = 32'h3c021040;
30'h00000014: inst = 32'h8fa30024;
30'h00000015: inst = 32'h00000000;
30'h00000016: inst = 32'h8fa40020;
30'h00000017: inst = 32'h00000000;
30'h00000018: inst = 32'h00031880;
30'h00000019: inst = 32'h34420000;
30'h0000001a: inst = 32'h00621021;
30'h0000001b: inst = 32'hac440000;
30'h0000001c: inst = 32'h8fa20024;
30'h0000001d: inst = 32'h00000000;
30'h0000001e: inst = 32'h24420001;
30'h0000001f: inst = 32'hafa20024;
30'h00000020: inst = 32'h0800140c;
30'h00000021: inst = 32'h00000000;
30'h00000022: inst = 32'h24020000;
30'h00000023: inst = 32'h27bd0028;
30'h00000024: inst = 32'h03e00008;
30'h00000025: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
